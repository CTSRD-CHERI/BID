// 2018, Alexandre Joannou, University of Cambridge

package BID;

import BID_Core :: *;
import BID_Utils :: *;
import BID_SimUtils :: *;
import BID_Interface :: *;
import BID_Collections :: *;

export BID_Core :: *;
export BID_Utils :: *;
export BID_SimUtils :: *;
export BID_Interface :: *;
export BID_Collections :: *;

endpackage: BID
