import "BDPI" function Bit#(64) sysTime ();
